magic
tech sky130A
magscale 1 2
timestamp 1655825574
<< obsli1 >>
rect 1104 2159 298816 297585
<< obsm1 >>
rect 14 2128 298816 297616
<< metal2 >>
rect 16118 299200 16174 300000
rect 49606 299200 49662 300000
rect 83094 299200 83150 300000
rect 115938 299200 115994 300000
rect 149426 299200 149482 300000
rect 182914 299200 182970 300000
rect 216402 299200 216458 300000
rect 249890 299200 249946 300000
rect 283378 299200 283434 300000
rect 18 0 74 800
rect 32862 0 32918 800
rect 66350 0 66406 800
rect 99838 0 99894 800
rect 133326 0 133382 800
rect 166814 0 166870 800
rect 199658 0 199714 800
rect 233146 0 233202 800
rect 266634 0 266690 800
<< obsm2 >>
rect 20 299144 16062 299200
rect 16230 299144 49550 299200
rect 49718 299144 83038 299200
rect 83206 299144 115882 299200
rect 116050 299144 149370 299200
rect 149538 299144 182858 299200
rect 183026 299144 216346 299200
rect 216514 299144 249834 299200
rect 250002 299144 283322 299200
rect 283490 299144 298154 299200
rect 20 856 298154 299144
rect 130 31 32806 856
rect 32974 31 66294 856
rect 66462 31 99782 856
rect 99950 31 133270 856
rect 133438 31 166758 856
rect 166926 31 199602 856
rect 199770 31 233090 856
rect 233258 31 266578 856
rect 266746 31 298154 856
<< metal3 >>
rect 299200 282208 300000 282328
rect 0 281528 800 281648
rect 299200 246848 300000 246968
rect 0 246168 800 246288
rect 299200 211488 300000 211608
rect 0 210808 800 210928
rect 0 176128 800 176248
rect 299200 176128 300000 176248
rect 0 140768 800 140888
rect 299200 140768 300000 140888
rect 0 105408 800 105528
rect 299200 105408 300000 105528
rect 299200 70728 300000 70848
rect 0 70048 800 70168
rect 299200 35368 300000 35488
rect 0 34688 800 34808
rect 299200 8 300000 128
<< obsm3 >>
rect 800 282408 299200 297601
rect 800 282128 299120 282408
rect 800 281728 299200 282128
rect 880 281448 299200 281728
rect 800 247048 299200 281448
rect 800 246768 299120 247048
rect 800 246368 299200 246768
rect 880 246088 299200 246368
rect 800 211688 299200 246088
rect 800 211408 299120 211688
rect 800 211008 299200 211408
rect 880 210728 299200 211008
rect 800 176328 299200 210728
rect 880 176048 299120 176328
rect 800 140968 299200 176048
rect 880 140688 299120 140968
rect 800 105608 299200 140688
rect 880 105328 299120 105608
rect 800 70928 299200 105328
rect 800 70648 299120 70928
rect 800 70248 299200 70648
rect 880 69968 299200 70248
rect 800 35568 299200 69968
rect 800 35288 299120 35568
rect 800 34888 299200 35288
rect 880 34608 299200 34888
rect 800 208 299200 34608
rect 800 35 299120 208
<< metal4 >>
rect 4208 2128 4528 297616
rect 19568 2128 19888 297616
rect 34928 2128 35248 297616
rect 50288 2128 50608 297616
rect 65648 2128 65968 297616
rect 81008 2128 81328 297616
rect 96368 2128 96688 297616
rect 111728 2128 112048 297616
rect 127088 2128 127408 297616
rect 142448 2128 142768 297616
rect 157808 2128 158128 297616
rect 173168 2128 173488 297616
rect 188528 2128 188848 297616
rect 203888 2128 204208 297616
rect 219248 2128 219568 297616
rect 234608 2128 234928 297616
rect 249968 2128 250288 297616
rect 265328 2128 265648 297616
rect 280688 2128 281008 297616
rect 296048 2128 296368 297616
<< obsm4 >>
rect 80835 6155 80928 297261
rect 81408 6155 96288 297261
rect 96768 6155 111648 297261
rect 112128 6155 127008 297261
rect 127488 6155 142368 297261
rect 142848 6155 157728 297261
rect 158208 6155 173088 297261
rect 173568 6155 188448 297261
rect 188928 6155 203808 297261
rect 204288 6155 219168 297261
rect 219648 6155 230861 297261
<< labels >>
rlabel metal2 s 83094 299200 83150 300000 6 address_bus[0]
port 1 nsew signal input
rlabel metal2 s 249890 299200 249946 300000 6 address_bus[1]
port 2 nsew signal input
rlabel metal2 s 16118 299200 16174 300000 6 address_bus[2]
port 3 nsew signal input
rlabel metal3 s 0 246168 800 246288 6 address_bus[3]
port 4 nsew signal input
rlabel metal2 s 233146 0 233202 800 6 address_bus[4]
port 5 nsew signal input
rlabel metal3 s 0 105408 800 105528 6 address_bus[5]
port 6 nsew signal input
rlabel metal2 s 216402 299200 216458 300000 6 address_bus[6]
port 7 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 address_bus[7]
port 8 nsew signal input
rlabel metal3 s 0 176128 800 176248 6 clk
port 9 nsew signal input
rlabel metal3 s 299200 211488 300000 211608 6 data_bus[0]
port 10 nsew signal input
rlabel metal3 s 299200 8 300000 128 6 data_bus[1]
port 11 nsew signal input
rlabel metal2 s 266634 0 266690 800 6 data_bus[2]
port 12 nsew signal input
rlabel metal3 s 0 70048 800 70168 6 data_bus[3]
port 13 nsew signal input
rlabel metal3 s 299200 176128 300000 176248 6 data_bus[4]
port 14 nsew signal input
rlabel metal2 s 18 0 74 800 6 data_bus[5]
port 15 nsew signal input
rlabel metal2 s 182914 299200 182970 300000 6 data_bus[6]
port 16 nsew signal input
rlabel metal3 s 299200 105408 300000 105528 6 data_bus[7]
port 17 nsew signal input
rlabel metal3 s 0 210808 800 210928 6 ext_write
port 18 nsew signal input
rlabel metal2 s 49606 299200 49662 300000 6 io_oeb[0]
port 19 nsew signal output
rlabel metal2 s 199658 0 199714 800 6 io_oeb[1]
port 20 nsew signal output
rlabel metal2 s 283378 299200 283434 300000 6 io_oeb[2]
port 21 nsew signal output
rlabel metal3 s 299200 35368 300000 35488 6 io_oeb[3]
port 22 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 io_oeb[4]
port 23 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 io_oeb[5]
port 24 nsew signal output
rlabel metal2 s 99838 0 99894 800 6 io_oeb[6]
port 25 nsew signal output
rlabel metal3 s 299200 70728 300000 70848 6 io_oeb[7]
port 26 nsew signal output
rlabel metal2 s 133326 0 133382 800 6 memory_bus[0]
port 27 nsew signal output
rlabel metal3 s 299200 246848 300000 246968 6 memory_bus[1]
port 28 nsew signal output
rlabel metal3 s 299200 282208 300000 282328 6 memory_bus[2]
port 29 nsew signal output
rlabel metal2 s 115938 299200 115994 300000 6 memory_bus[3]
port 30 nsew signal output
rlabel metal2 s 149426 299200 149482 300000 6 memory_bus[4]
port 31 nsew signal output
rlabel metal2 s 166814 0 166870 800 6 memory_bus[5]
port 32 nsew signal output
rlabel metal3 s 0 140768 800 140888 6 memory_bus[6]
port 33 nsew signal output
rlabel metal3 s 0 281528 800 281648 6 memory_bus[7]
port 34 nsew signal output
rlabel metal3 s 299200 140768 300000 140888 6 rst
port 35 nsew signal input
rlabel metal4 s 4208 2128 4528 297616 6 vccd1
port 36 nsew power input
rlabel metal4 s 34928 2128 35248 297616 6 vccd1
port 36 nsew power input
rlabel metal4 s 65648 2128 65968 297616 6 vccd1
port 36 nsew power input
rlabel metal4 s 96368 2128 96688 297616 6 vccd1
port 36 nsew power input
rlabel metal4 s 127088 2128 127408 297616 6 vccd1
port 36 nsew power input
rlabel metal4 s 157808 2128 158128 297616 6 vccd1
port 36 nsew power input
rlabel metal4 s 188528 2128 188848 297616 6 vccd1
port 36 nsew power input
rlabel metal4 s 219248 2128 219568 297616 6 vccd1
port 36 nsew power input
rlabel metal4 s 249968 2128 250288 297616 6 vccd1
port 36 nsew power input
rlabel metal4 s 280688 2128 281008 297616 6 vccd1
port 36 nsew power input
rlabel metal4 s 19568 2128 19888 297616 6 vssd1
port 37 nsew ground input
rlabel metal4 s 50288 2128 50608 297616 6 vssd1
port 37 nsew ground input
rlabel metal4 s 81008 2128 81328 297616 6 vssd1
port 37 nsew ground input
rlabel metal4 s 111728 2128 112048 297616 6 vssd1
port 37 nsew ground input
rlabel metal4 s 142448 2128 142768 297616 6 vssd1
port 37 nsew ground input
rlabel metal4 s 173168 2128 173488 297616 6 vssd1
port 37 nsew ground input
rlabel metal4 s 203888 2128 204208 297616 6 vssd1
port 37 nsew ground input
rlabel metal4 s 234608 2128 234928 297616 6 vssd1
port 37 nsew ground input
rlabel metal4 s 265328 2128 265648 297616 6 vssd1
port 37 nsew ground input
rlabel metal4 s 296048 2128 296368 297616 6 vssd1
port 37 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 300000 300000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 68568574
string GDS_FILE /home/mdtanvirarafin/caravel_user_project/openlane/risc_spm/runs/risc_spm/results/finishing/RISC_SPM.magic.gds
string GDS_START 1100726
<< end >>

