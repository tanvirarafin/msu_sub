VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RISC_SPM
  CLASS BLOCK ;
  FOREIGN RISC_SPM ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 1500.000 ;
  PIN address_bus[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 1496.000 415.750 1500.000 ;
    END
  END address_bus[0]
  PIN address_bus[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.450 1496.000 1249.730 1500.000 ;
    END
  END address_bus[1]
  PIN address_bus[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 1496.000 80.870 1500.000 ;
    END
  END address_bus[2]
  PIN address_bus[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1230.840 4.000 1231.440 ;
    END
  END address_bus[3]
  PIN address_bus[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.730 0.000 1166.010 4.000 ;
    END
  END address_bus[4]
  PIN address_bus[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.040 4.000 527.640 ;
    END
  END address_bus[5]
  PIN address_bus[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.010 1496.000 1082.290 1500.000 ;
    END
  END address_bus[6]
  PIN address_bus[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END address_bus[7]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 880.640 4.000 881.240 ;
    END
  END clk
  PIN data_bus[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1057.440 1500.000 1058.040 ;
    END
  END data_bus[0]
  PIN data_bus[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 0.040 1500.000 0.640 ;
    END
  END data_bus[1]
  PIN data_bus[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.170 0.000 1333.450 4.000 ;
    END
  END data_bus[2]
  PIN data_bus[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END data_bus[3]
  PIN data_bus[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 880.640 1500.000 881.240 ;
    END
  END data_bus[4]
  PIN data_bus[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END data_bus[5]
  PIN data_bus[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.570 1496.000 914.850 1500.000 ;
    END
  END data_bus[6]
  PIN data_bus[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 527.040 1500.000 527.640 ;
    END
  END data_bus[7]
  PIN ext_write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1054.040 4.000 1054.640 ;
    END
  END ext_write
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 1496.000 248.310 1500.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.290 0.000 998.570 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1416.890 1496.000 1417.170 1500.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 176.840 1500.000 177.440 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 0.000 499.470 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 353.640 1500.000 354.240 ;
    END
  END io_oeb[7]
  PIN memory_bus[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 0.000 666.910 4.000 ;
    END
  END memory_bus[0]
  PIN memory_bus[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1234.240 1500.000 1234.840 ;
    END
  END memory_bus[1]
  PIN memory_bus[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1411.040 1500.000 1411.640 ;
    END
  END memory_bus[2]
  PIN memory_bus[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 1496.000 579.970 1500.000 ;
    END
  END memory_bus[3]
  PIN memory_bus[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 1496.000 747.410 1500.000 ;
    END
  END memory_bus[4]
  PIN memory_bus[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.070 0.000 834.350 4.000 ;
    END
  END memory_bus[5]
  PIN memory_bus[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.840 4.000 704.440 ;
    END
  END memory_bus[6]
  PIN memory_bus[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1407.640 4.000 1408.240 ;
    END
  END memory_bus[7]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 703.840 1500.000 704.440 ;
    END
  END rst
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1488.080 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1494.080 1487.925 ;
      LAYER met1 ;
        RECT 0.070 10.640 1494.080 1488.080 ;
      LAYER met2 ;
        RECT 0.100 1495.720 80.310 1496.000 ;
        RECT 81.150 1495.720 247.750 1496.000 ;
        RECT 248.590 1495.720 415.190 1496.000 ;
        RECT 416.030 1495.720 579.410 1496.000 ;
        RECT 580.250 1495.720 746.850 1496.000 ;
        RECT 747.690 1495.720 914.290 1496.000 ;
        RECT 915.130 1495.720 1081.730 1496.000 ;
        RECT 1082.570 1495.720 1249.170 1496.000 ;
        RECT 1250.010 1495.720 1416.610 1496.000 ;
        RECT 1417.450 1495.720 1490.770 1496.000 ;
        RECT 0.100 4.280 1490.770 1495.720 ;
        RECT 0.650 0.155 164.030 4.280 ;
        RECT 164.870 0.155 331.470 4.280 ;
        RECT 332.310 0.155 498.910 4.280 ;
        RECT 499.750 0.155 666.350 4.280 ;
        RECT 667.190 0.155 833.790 4.280 ;
        RECT 834.630 0.155 998.010 4.280 ;
        RECT 998.850 0.155 1165.450 4.280 ;
        RECT 1166.290 0.155 1332.890 4.280 ;
        RECT 1333.730 0.155 1490.770 4.280 ;
      LAYER met3 ;
        RECT 4.000 1412.040 1496.000 1488.005 ;
        RECT 4.000 1410.640 1495.600 1412.040 ;
        RECT 4.000 1408.640 1496.000 1410.640 ;
        RECT 4.400 1407.240 1496.000 1408.640 ;
        RECT 4.000 1235.240 1496.000 1407.240 ;
        RECT 4.000 1233.840 1495.600 1235.240 ;
        RECT 4.000 1231.840 1496.000 1233.840 ;
        RECT 4.400 1230.440 1496.000 1231.840 ;
        RECT 4.000 1058.440 1496.000 1230.440 ;
        RECT 4.000 1057.040 1495.600 1058.440 ;
        RECT 4.000 1055.040 1496.000 1057.040 ;
        RECT 4.400 1053.640 1496.000 1055.040 ;
        RECT 4.000 881.640 1496.000 1053.640 ;
        RECT 4.400 880.240 1495.600 881.640 ;
        RECT 4.000 704.840 1496.000 880.240 ;
        RECT 4.400 703.440 1495.600 704.840 ;
        RECT 4.000 528.040 1496.000 703.440 ;
        RECT 4.400 526.640 1495.600 528.040 ;
        RECT 4.000 354.640 1496.000 526.640 ;
        RECT 4.000 353.240 1495.600 354.640 ;
        RECT 4.000 351.240 1496.000 353.240 ;
        RECT 4.400 349.840 1496.000 351.240 ;
        RECT 4.000 177.840 1496.000 349.840 ;
        RECT 4.000 176.440 1495.600 177.840 ;
        RECT 4.000 174.440 1496.000 176.440 ;
        RECT 4.400 173.040 1496.000 174.440 ;
        RECT 4.000 1.040 1496.000 173.040 ;
        RECT 4.000 0.175 1495.600 1.040 ;
      LAYER met4 ;
        RECT 419.815 11.735 481.440 1486.305 ;
        RECT 483.840 11.735 558.240 1486.305 ;
        RECT 560.640 11.735 635.040 1486.305 ;
        RECT 637.440 11.735 711.840 1486.305 ;
        RECT 714.240 11.735 788.640 1486.305 ;
        RECT 791.040 11.735 865.440 1486.305 ;
        RECT 867.840 11.735 942.240 1486.305 ;
        RECT 944.640 11.735 1019.040 1486.305 ;
        RECT 1021.440 11.735 1095.840 1486.305 ;
        RECT 1098.240 11.735 1126.705 1486.305 ;
  END
END RISC_SPM
END LIBRARY

