VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RISC_SPM
  CLASS BLOCK ;
  FOREIGN RISC_SPM ;
  ORIGIN 0.000 0.000 ;
  SIZE 1000.000 BY 1000.000 ;
  PIN address_bus[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 996.000 277.290 1000.000 ;
    END
  END address_bus[0]
  PIN address_bus[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.070 996.000 834.350 1000.000 ;
    END
  END address_bus[1]
  PIN address_bus[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 996.000 55.110 1000.000 ;
    END
  END address_bus[2]
  PIN address_bus[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 819.440 4.000 820.040 ;
    END
  END address_bus[3]
  PIN address_bus[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 0.000 779.610 4.000 ;
    END
  END address_bus[4]
  PIN address_bus[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END address_bus[5]
  PIN address_bus[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 996.000 721.650 1000.000 ;
    END
  END address_bus[6]
  PIN address_bus[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END address_bus[7]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END clk
  PIN data_bus[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 703.840 1000.000 704.440 ;
    END
  END data_bus[0]
  PIN data_bus[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 0.040 1000.000 0.640 ;
    END
  END data_bus[1]
  PIN data_bus[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 0.000 889.090 4.000 ;
    END
  END data_bus[2]
  PIN data_bus[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END data_bus[3]
  PIN data_bus[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 588.240 1000.000 588.840 ;
    END
  END data_bus[4]
  PIN data_bus[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END data_bus[5]
  PIN data_bus[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 996.000 608.950 1000.000 ;
    END
  END data_bus[6]
  PIN data_bus[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 350.240 1000.000 350.840 ;
    END
  END data_bus[7]
  PIN ext_write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.840 4.000 704.440 ;
    END
  END ext_write
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 996.000 164.590 1000.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 0.000 666.910 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 996.000 943.830 1000.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 115.640 1000.000 116.240 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 234.640 1000.000 235.240 ;
    END
  END io_oeb[7]
  PIN memory_bus[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END memory_bus[0]
  PIN memory_bus[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 822.840 1000.000 823.440 ;
    END
  END memory_bus[1]
  PIN memory_bus[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 938.440 1000.000 939.040 ;
    END
  END memory_bus[2]
  PIN memory_bus[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 996.000 386.770 1000.000 ;
    END
  END memory_bus[3]
  PIN memory_bus[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 996.000 499.470 1000.000 ;
    END
  END memory_bus[4]
  PIN memory_bus[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 0.000 554.210 4.000 ;
    END
  END memory_bus[5]
  PIN memory_bus[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END memory_bus[6]
  PIN memory_bus[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 938.440 4.000 939.040 ;
    END
  END memory_bus[7]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 469.240 1000.000 469.840 ;
    END
  END rst
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 987.600 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 987.600 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 994.060 987.445 ;
      LAYER met1 ;
        RECT 0.070 10.640 994.060 987.600 ;
      LAYER met2 ;
        RECT 0.100 995.720 54.550 996.610 ;
        RECT 55.390 995.720 164.030 996.610 ;
        RECT 164.870 995.720 276.730 996.610 ;
        RECT 277.570 995.720 386.210 996.610 ;
        RECT 387.050 995.720 498.910 996.610 ;
        RECT 499.750 995.720 608.390 996.610 ;
        RECT 609.230 995.720 721.090 996.610 ;
        RECT 721.930 995.720 833.790 996.610 ;
        RECT 834.630 995.720 943.270 996.610 ;
        RECT 944.110 995.720 990.750 996.610 ;
        RECT 0.100 4.280 990.750 995.720 ;
        RECT 0.650 0.155 109.290 4.280 ;
        RECT 110.130 0.155 221.990 4.280 ;
        RECT 222.830 0.155 331.470 4.280 ;
        RECT 332.310 0.155 444.170 4.280 ;
        RECT 445.010 0.155 553.650 4.280 ;
        RECT 554.490 0.155 666.350 4.280 ;
        RECT 667.190 0.155 779.050 4.280 ;
        RECT 779.890 0.155 888.530 4.280 ;
        RECT 889.370 0.155 990.750 4.280 ;
      LAYER met3 ;
        RECT 4.000 939.440 996.000 987.525 ;
        RECT 4.400 938.040 995.600 939.440 ;
        RECT 4.000 823.840 996.000 938.040 ;
        RECT 4.000 822.440 995.600 823.840 ;
        RECT 4.000 820.440 996.000 822.440 ;
        RECT 4.400 819.040 996.000 820.440 ;
        RECT 4.000 704.840 996.000 819.040 ;
        RECT 4.400 703.440 995.600 704.840 ;
        RECT 4.000 589.240 996.000 703.440 ;
        RECT 4.000 587.840 995.600 589.240 ;
        RECT 4.000 585.840 996.000 587.840 ;
        RECT 4.400 584.440 996.000 585.840 ;
        RECT 4.000 470.240 996.000 584.440 ;
        RECT 4.400 468.840 995.600 470.240 ;
        RECT 4.000 351.240 996.000 468.840 ;
        RECT 4.400 349.840 995.600 351.240 ;
        RECT 4.000 235.640 996.000 349.840 ;
        RECT 4.400 234.240 995.600 235.640 ;
        RECT 4.000 116.640 996.000 234.240 ;
        RECT 4.400 115.240 995.600 116.640 ;
        RECT 4.000 1.040 996.000 115.240 ;
        RECT 4.000 0.175 995.600 1.040 ;
      LAYER met4 ;
        RECT 86.775 11.735 97.440 985.825 ;
        RECT 99.840 11.735 174.240 985.825 ;
        RECT 176.640 11.735 251.040 985.825 ;
        RECT 253.440 11.735 327.840 985.825 ;
        RECT 330.240 11.735 404.640 985.825 ;
        RECT 407.040 11.735 481.440 985.825 ;
        RECT 483.840 11.735 558.240 985.825 ;
        RECT 560.640 11.735 635.040 985.825 ;
        RECT 637.440 11.735 711.840 985.825 ;
        RECT 714.240 11.735 784.465 985.825 ;
  END
END RISC_SPM
END LIBRARY

