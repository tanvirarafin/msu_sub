VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO asmd_multiplier
  CLASS BLOCK ;
  FOREIGN asmd_multiplier ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 51.040 300.000 51.640 ;
    END
  END clk
  PIN product[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 296.000 299.830 300.000 ;
    END
  END product[0]
  PIN product[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 296.000 183.910 300.000 ;
    END
  END product[1]
  PIN product[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END product[2]
  PIN product[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 238.040 300.000 238.640 ;
    END
  END product[3]
  PIN product[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END product[4]
  PIN product[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END product[5]
  PIN product[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 296.000 125.950 300.000 ;
    END
  END product[6]
  PIN product[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END product[7]
  PIN ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 296.000 64.770 300.000 ;
    END
  END ready
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END reset
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END start
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
  END vssd1
  PIN word0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END word0[0]
  PIN word0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 176.840 300.000 177.440 ;
    END
  END word0[1]
  PIN word0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END word0[2]
  PIN word0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 296.000 241.870 300.000 ;
    END
  END word0[3]
  PIN word1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END word1[0]
  PIN word1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END word1[1]
  PIN word1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 296.000 6.810 300.000 ;
    END
  END word1[2]
  PIN word1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 115.640 300.000 116.240 ;
    END
  END word1[3]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 294.400 288.405 ;
      LAYER met1 ;
        RECT 0.070 10.640 299.850 288.560 ;
      LAYER met2 ;
        RECT 0.100 295.720 6.250 296.210 ;
        RECT 7.090 295.720 64.210 296.210 ;
        RECT 65.050 295.720 125.390 296.210 ;
        RECT 126.230 295.720 183.350 296.210 ;
        RECT 184.190 295.720 241.310 296.210 ;
        RECT 242.150 295.720 299.270 296.210 ;
        RECT 0.100 4.280 299.820 295.720 ;
        RECT 0.650 4.000 57.770 4.280 ;
        RECT 58.610 4.000 115.730 4.280 ;
        RECT 116.570 4.000 173.690 4.280 ;
        RECT 174.530 4.000 234.870 4.280 ;
        RECT 235.710 4.000 292.830 4.280 ;
        RECT 293.670 4.000 299.820 4.280 ;
      LAYER met3 ;
        RECT 4.000 249.240 296.000 288.485 ;
        RECT 4.400 247.840 296.000 249.240 ;
        RECT 4.000 239.040 296.000 247.840 ;
        RECT 4.000 237.640 295.600 239.040 ;
        RECT 4.000 184.640 296.000 237.640 ;
        RECT 4.400 183.240 296.000 184.640 ;
        RECT 4.000 177.840 296.000 183.240 ;
        RECT 4.000 176.440 295.600 177.840 ;
        RECT 4.000 123.440 296.000 176.440 ;
        RECT 4.400 122.040 296.000 123.440 ;
        RECT 4.000 116.640 296.000 122.040 ;
        RECT 4.000 115.240 295.600 116.640 ;
        RECT 4.000 62.240 296.000 115.240 ;
        RECT 4.400 60.840 296.000 62.240 ;
        RECT 4.000 52.040 296.000 60.840 ;
        RECT 4.000 50.640 295.600 52.040 ;
        RECT 4.000 10.715 296.000 50.640 ;
  END
END asmd_multiplier
END LIBRARY

