magic
tech sky130A
timestamp 1608324878
<< checkpaint >>
rect 1495 5490 6500 6570
rect -630 428 19262 5490
rect -630 -630 6210 428
rect 16092 356 18972 428
<< fillblock >>
rect -328 754 16860 5172
use alpha_D  alphaX_0 hexdigits
timestamp 1598786981
transform 1 0 14887 0 1 1080
box 0 0 1620 3780
use alpha_C  alphaX_1 hexdigits
timestamp 1598786981
transform 1 0 12750 0 1 1080
box 0 0 1620 3780
use alpha_B  alphaX_2 hexdigits
timestamp 1598786981
transform 1 0 10625 0 1 1080
box 0 0 1620 3780
use alpha_A  alphaX_3 hexdigits
timestamp 1598786981
transform 1 0 8500 0 1 1080
box 0 0 1620 3780
use alpha_0  alphaX_4 hexdigits
timestamp 1598786981
transform 1 0 6375 0 1 1080
box 0 0 1620 3780
use alpha_0  alphaX_5
timestamp 1598786981
transform 1 0 4250 0 1 1080
box 0 0 1620 3780
use alpha_0  alphaX_6
timestamp 1598786981
transform 1 0 2125 0 1 1080
box 0 0 1620 3780
use alpha_0  alphaX_7
timestamp 1598786981
transform 1 0 0 0 1 1080
box 0 0 1620 3780
<< end >>
