magic
tech sky130A
magscale 1 2
timestamp 1655863783
<< obsli1 >>
rect 1104 2159 198812 197489
<< obsm1 >>
rect 14 2128 198812 197520
<< metal2 >>
rect 10966 199200 11022 200000
rect 32862 199200 32918 200000
rect 55402 199200 55458 200000
rect 77298 199200 77354 200000
rect 99838 199200 99894 200000
rect 121734 199200 121790 200000
rect 144274 199200 144330 200000
rect 166814 199200 166870 200000
rect 188710 199200 188766 200000
rect 18 0 74 800
rect 21914 0 21970 800
rect 44454 0 44510 800
rect 66350 0 66406 800
rect 88890 0 88946 800
rect 110786 0 110842 800
rect 133326 0 133382 800
rect 155866 0 155922 800
rect 177762 0 177818 800
<< obsm2 >>
rect 20 199144 10910 199322
rect 11078 199144 32806 199322
rect 32974 199144 55346 199322
rect 55514 199144 77242 199322
rect 77410 199144 99782 199322
rect 99950 199144 121678 199322
rect 121846 199144 144218 199322
rect 144386 199144 166758 199322
rect 166926 199144 188654 199322
rect 188822 199144 198150 199322
rect 20 856 198150 199144
rect 130 31 21858 856
rect 22026 31 44398 856
rect 44566 31 66294 856
rect 66462 31 88834 856
rect 89002 31 110730 856
rect 110898 31 133270 856
rect 133438 31 155810 856
rect 155978 31 177706 856
rect 177874 31 198150 856
<< metal3 >>
rect 0 187688 800 187808
rect 199200 187688 200000 187808
rect 199200 164568 200000 164688
rect 0 163888 800 164008
rect 0 140768 800 140888
rect 199200 140768 200000 140888
rect 199200 117648 200000 117768
rect 0 116968 800 117088
rect 0 93848 800 93968
rect 199200 93848 200000 93968
rect 0 70048 800 70168
rect 199200 70048 200000 70168
rect 0 46928 800 47048
rect 199200 46928 200000 47048
rect 0 23128 800 23248
rect 199200 23128 200000 23248
rect 199200 8 200000 128
<< obsm3 >>
rect 800 187888 199200 197505
rect 880 187608 199120 187888
rect 800 164768 199200 187608
rect 800 164488 199120 164768
rect 800 164088 199200 164488
rect 880 163808 199200 164088
rect 800 140968 199200 163808
rect 880 140688 199120 140968
rect 800 117848 199200 140688
rect 800 117568 199120 117848
rect 800 117168 199200 117568
rect 880 116888 199200 117168
rect 800 94048 199200 116888
rect 880 93768 199120 94048
rect 800 70248 199200 93768
rect 880 69968 199120 70248
rect 800 47128 199200 69968
rect 880 46848 199120 47128
rect 800 23328 199200 46848
rect 880 23048 199120 23328
rect 800 208 199200 23048
rect 800 35 199120 208
<< metal4 >>
rect 4208 2128 4528 197520
rect 19568 2128 19888 197520
rect 34928 2128 35248 197520
rect 50288 2128 50608 197520
rect 65648 2128 65968 197520
rect 81008 2128 81328 197520
rect 96368 2128 96688 197520
rect 111728 2128 112048 197520
rect 127088 2128 127408 197520
rect 142448 2128 142768 197520
rect 157808 2128 158128 197520
rect 173168 2128 173488 197520
rect 188528 2128 188848 197520
<< obsm4 >>
rect 17355 2347 19488 197165
rect 19968 2347 34848 197165
rect 35328 2347 50208 197165
rect 50688 2347 65568 197165
rect 66048 2347 80928 197165
rect 81408 2347 96288 197165
rect 96768 2347 111648 197165
rect 112128 2347 127008 197165
rect 127488 2347 142368 197165
rect 142848 2347 156893 197165
<< labels >>
rlabel metal2 s 55402 199200 55458 200000 6 address_bus[0]
port 1 nsew signal input
rlabel metal2 s 166814 199200 166870 200000 6 address_bus[1]
port 2 nsew signal input
rlabel metal2 s 10966 199200 11022 200000 6 address_bus[2]
port 3 nsew signal input
rlabel metal3 s 0 163888 800 164008 6 address_bus[3]
port 4 nsew signal input
rlabel metal2 s 155866 0 155922 800 6 address_bus[4]
port 5 nsew signal input
rlabel metal3 s 0 70048 800 70168 6 address_bus[5]
port 6 nsew signal input
rlabel metal2 s 144274 199200 144330 200000 6 address_bus[6]
port 7 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 address_bus[7]
port 8 nsew signal input
rlabel metal3 s 0 116968 800 117088 6 clk
port 9 nsew signal input
rlabel metal3 s 199200 140768 200000 140888 6 data_bus[0]
port 10 nsew signal input
rlabel metal3 s 199200 8 200000 128 6 data_bus[1]
port 11 nsew signal input
rlabel metal2 s 177762 0 177818 800 6 data_bus[2]
port 12 nsew signal input
rlabel metal3 s 0 46928 800 47048 6 data_bus[3]
port 13 nsew signal input
rlabel metal3 s 199200 117648 200000 117768 6 data_bus[4]
port 14 nsew signal input
rlabel metal2 s 18 0 74 800 6 data_bus[5]
port 15 nsew signal input
rlabel metal2 s 121734 199200 121790 200000 6 data_bus[6]
port 16 nsew signal input
rlabel metal3 s 199200 70048 200000 70168 6 data_bus[7]
port 17 nsew signal input
rlabel metal3 s 0 140768 800 140888 6 ext_write
port 18 nsew signal input
rlabel metal2 s 32862 199200 32918 200000 6 io_oeb[0]
port 19 nsew signal output
rlabel metal2 s 133326 0 133382 800 6 io_oeb[1]
port 20 nsew signal output
rlabel metal2 s 188710 199200 188766 200000 6 io_oeb[2]
port 21 nsew signal output
rlabel metal3 s 199200 23128 200000 23248 6 io_oeb[3]
port 22 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 io_oeb[4]
port 23 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 io_oeb[5]
port 24 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 io_oeb[6]
port 25 nsew signal output
rlabel metal3 s 199200 46928 200000 47048 6 io_oeb[7]
port 26 nsew signal output
rlabel metal2 s 88890 0 88946 800 6 memory_bus[0]
port 27 nsew signal output
rlabel metal3 s 199200 164568 200000 164688 6 memory_bus[1]
port 28 nsew signal output
rlabel metal3 s 199200 187688 200000 187808 6 memory_bus[2]
port 29 nsew signal output
rlabel metal2 s 77298 199200 77354 200000 6 memory_bus[3]
port 30 nsew signal output
rlabel metal2 s 99838 199200 99894 200000 6 memory_bus[4]
port 31 nsew signal output
rlabel metal2 s 110786 0 110842 800 6 memory_bus[5]
port 32 nsew signal output
rlabel metal3 s 0 93848 800 93968 6 memory_bus[6]
port 33 nsew signal output
rlabel metal3 s 0 187688 800 187808 6 memory_bus[7]
port 34 nsew signal output
rlabel metal3 s 199200 93848 200000 93968 6 rst
port 35 nsew signal input
rlabel metal4 s 4208 2128 4528 197520 6 vccd1
port 36 nsew power input
rlabel metal4 s 34928 2128 35248 197520 6 vccd1
port 36 nsew power input
rlabel metal4 s 65648 2128 65968 197520 6 vccd1
port 36 nsew power input
rlabel metal4 s 96368 2128 96688 197520 6 vccd1
port 36 nsew power input
rlabel metal4 s 127088 2128 127408 197520 6 vccd1
port 36 nsew power input
rlabel metal4 s 157808 2128 158128 197520 6 vccd1
port 36 nsew power input
rlabel metal4 s 188528 2128 188848 197520 6 vccd1
port 36 nsew power input
rlabel metal4 s 19568 2128 19888 197520 6 vssd1
port 37 nsew ground input
rlabel metal4 s 50288 2128 50608 197520 6 vssd1
port 37 nsew ground input
rlabel metal4 s 81008 2128 81328 197520 6 vssd1
port 37 nsew ground input
rlabel metal4 s 111728 2128 112048 197520 6 vssd1
port 37 nsew ground input
rlabel metal4 s 142448 2128 142768 197520 6 vssd1
port 37 nsew ground input
rlabel metal4 s 173168 2128 173488 197520 6 vssd1
port 37 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 200000 200000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 56239092
string GDS_FILE /home/mdtanvirarafin/caravel_user_project/openlane/risc_spm/runs/risc_spm/results/finishing/RISC_SPM.magic.gds
string GDS_START 1075618
<< end >>

